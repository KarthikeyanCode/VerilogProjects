//have to work on this
module serial_adder();